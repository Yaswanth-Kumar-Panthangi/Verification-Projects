package bridge_pkg;

     import uvm_pkg::*;
	 `include "uvm_macros.svh"
	 
	 `include "ahb_config.sv"
	 `include "apb_config.sv"
	 `include "env_config.sv"
	 
	 `include "ahb_xtn.sv"
     	 `include "ahb_seq.sv"
	 `include "ahb_sequencer.sv"
	 `include "ahb_driver.sv"
	 `include "ahb_monitor.sv"
	 `include "ahb_agt.sv"
	 `include "ahb_agt_top.sv"
	 
	 `include "apb_xtn.sv"
	 `include "apb_sequencer.sv"
	 `include "apb_driver.sv"
	 `include "apb_monitor.sv"
	 `include "apb_agt.sv"
	 `include "apb_agt_top.sv"
	 `include "sb.sv"
	 `include "env.sv"
	 `include "test.sv"
endpackage
